module vga3_top(
    input r,
    input g,
    input b,
    input hsync,
    input vsync
);

    

endmodule



