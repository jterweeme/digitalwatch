module buttons(
    input csi_clk,
    input csi_rst,
);

endmodule


