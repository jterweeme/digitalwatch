library ieee;
use ieee.std_logic_1164.all;

entity myrtc is
    port (clk, reset: in std_logic);
end myrtc;

architecture behavior of myrtc is
begin
    
end behavior;


